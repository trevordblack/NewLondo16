module loadhex();




endmodule