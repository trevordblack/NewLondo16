module fetch(C, A, B, loadHex, 3op, valueC, valueA, valueB);
	input [3:0] C, A, B;
	input loadHex, 3op;
	output [31:0] valueC, valueA, valueB;
	output [2:0] request
	
	
endmodule