module newlondo();
	
	instruction_fetch();
	decode();
	register_fetch();
	execute();
	write_back();
	
endmodule